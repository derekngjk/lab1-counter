module counter # (
    parameter WIDTH = 8
) (
    // interface signals
    input logic             clk,
    input logic             rst,
    input logic             en,
    output logic[WIDTH-1:0] count
);

/*
Default implementation: if rst is high set count to 0
Else increment count by en
*/
always_ff @ (posedge clk)
    if (rst) count <= {WIDTH{1'b0}};
    else     count <= count + {{WIDTH-1{1'b0}}, en};


endmodule
